CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 963
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 114 299 0 1 11
0 8
0
0 0 20592 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
43551.5 0
0
13 Logic Switch~
5 114 265 0 1 11
0 7
0
0 0 20592 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3472 0 0
2
43551.5 0
0
14 Logic Display~
6 714 257 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
6 SumOut
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
43551.5 0
0
14 Logic Display~
6 662 201 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
7 CarryOu
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3536 0 0
2
43551.5 0
0
5 4001~
219 538 275 0 3 22
0 3 4 2
0
0 0 624 0
4 4001
-14 -24 14 -16
5 Nor1A
-9 -25 26 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
4597 0 0
2
43551.5 0
0
5 4001~
219 448 236 0 3 22
0 6 5 3
0
0 0 624 0
4 4001
-14 -24 14 -16
4 NorD
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 1 0
1 U
3835 0 0
2
43551.5 1
0
5 4001~
219 274 376 0 3 22
0 8 8 5
0
0 0 624 0
4 4001
-14 -24 14 -16
4 NorC
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 1 0
1 U
3670 0 0
2
43551.5 0
0
5 4001~
219 278 286 0 3 22
0 7 8 4
0
0 0 624 0
4 4001
-14 -24 14 -16
4 NorB
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 1 0
1 U
5616 0 0
2
43551.5 0
0
5 4001~
219 275 205 0 3 22
0 7 7 6
0
0 0 624 0
4 4001
-14 -24 14 -16
4 NorA
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 1 0
1 U
9323 0 0
2
43551.5 0
0
12
3 1 2 0 0 4224 0 5 3 0 0 5
577 275
702 275
702 283
714 283
714 275
0 1 3 0 0 8320 0 0 4 4 0 4
517 236
517 227
662 227
662 219
3 2 4 0 0 4224 0 8 5 0 0 4
317 286
512 286
512 284
525 284
3 1 3 0 0 0 0 6 5 0 0 4
487 236
517 236
517 266
525 266
3 2 5 0 0 8320 0 7 6 0 0 4
313 376
427 376
427 245
435 245
3 1 6 0 0 4224 0 9 6 0 0 4
314 205
427 205
427 227
435 227
0 0 7 0 0 4096 0 0 0 12 9 3
228 265
228 202
254 202
0 0 8 0 0 4096 0 0 0 11 10 3
226 299
226 376
253 376
2 1 7 0 0 0 0 9 9 0 0 4
262 214
254 214
254 196
262 196
1 2 8 0 0 0 0 7 7 0 0 4
261 367
253 367
253 385
261 385
1 2 8 0 0 4224 0 1 8 0 0 4
126 299
257 299
257 295
265 295
1 1 7 0 0 4224 0 2 8 0 0 4
126 265
257 265
257 277
265 277
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
