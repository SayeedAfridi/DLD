CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 963
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 184 289 0 1 11
0 7
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3751 0 0
2
43551.5 0
0
13 Logic Switch~
5 181 246 0 1 11
0 8
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4292 0 0
2
43551.5 0
0
14 Logic Display~
6 826 250 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
7 DiffOut
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6118 0 0
2
43551.5 0
0
14 Logic Display~
6 615 173 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
6 Borrow
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
34 0 0
2
43551.5 0
0
5 4001~
219 712 273 0 3 22
0 4 4 2
0
0 0 624 0
4 4001
-14 -24 14 -16
5 Nor1A
-9 -25 26 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
6357 0 0
2
43551.5 0
0
5 4001~
219 470 340 0 3 22
0 6 7 5
0
0 0 624 0
4 4001
-14 -24 14 -16
4 NorD
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 1 0
1 U
319 0 0
2
43551.5 1
0
5 4001~
219 467 191 0 3 22
0 8 6 3
0
0 0 624 0
4 4001
-14 -24 14 -16
4 NorC
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 1 0
1 U
3976 0 0
2
43551.5 0
0
5 4001~
219 577 271 0 3 22
0 3 5 4
0
0 0 624 0
4 4001
-14 -24 14 -16
4 NorB
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 1 0
1 U
7634 0 0
2
43551.5 0
0
5 4001~
219 324 268 0 3 22
0 8 7 6
0
0 0 624 0
4 4001
-14 -24 14 -16
4 NorA
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 1 0
1 U
523 0 0
2
43551.5 0
0
12
1 3 2 0 0 8320 0 3 5 0 0 3
826 268
826 273
751 273
0 1 3 0 0 4224 0 0 4 5 0 2
514 191
615 191
3 0 4 0 0 4224 0 8 0 0 4 2
616 271
691 271
1 2 4 0 0 0 0 5 5 0 0 4
699 264
691 264
691 282
699 282
1 3 3 0 0 0 0 8 7 0 0 4
564 262
514 262
514 191
506 191
3 2 5 0 0 8320 0 6 8 0 0 4
509 340
556 340
556 280
564 280
3 0 6 0 0 4096 0 9 0 0 8 2
363 268
446 268
1 2 6 0 0 8320 0 6 7 0 0 4
457 331
446 331
446 200
454 200
0 2 7 0 0 8320 0 0 6 11 0 3
266 289
266 349
457 349
0 1 8 0 0 8320 0 0 7 12 0 3
266 246
266 182
454 182
1 2 7 0 0 0 0 1 9 0 0 4
196 289
303 289
303 277
311 277
1 1 8 0 0 0 0 2 9 0 0 4
193 246
303 246
303 259
311 259
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
