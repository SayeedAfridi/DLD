CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 963
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
6
13 Logic Switch~
5 197 261 0 1 11
0 5
0
0 0 20592 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
961 0 0
2
43551.5 0
0
13 Logic Switch~
5 196 206 0 1 11
0 4
0
0 0 20592 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3178 0 0
2
43551.5 0
0
14 Logic Display~
6 558 297 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
7 CarryOu
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3409 0 0
2
43551.5 0
0
14 Logic Display~
6 545 197 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
6 SumOut
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3951 0 0
2
43551.5 0
0
5 4081~
219 420 306 0 3 22
0 4 5 3
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
8885 0 0
2
43551.5 0
0
5 4030~
219 410 221 0 3 22
0 4 5 2
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3780 0 0
2
43551.5 0
0
6
3 1 2 0 0 4224 0 6 4 0 0 3
443 221
545 221
545 215
3 1 3 0 0 4224 0 5 3 0 0 5
441 306
546 306
546 323
558 323
558 315
0 1 4 0 0 8192 0 0 5 6 0 3
304 206
304 297
396 297
0 2 5 0 0 8192 0 0 5 5 0 3
252 261
252 315
396 315
1 2 5 0 0 4224 0 1 6 0 0 4
209 261
386 261
386 230
394 230
1 1 4 0 0 4224 0 2 6 0 0 4
208 206
386 206
386 212
394 212
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
