CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 963
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 149 247 0 1 11
0 6
0
0 0 21104 0
2 0V
-6 -16 8 -8
3 Cin
-13 -19 8 -11
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43551.5 0
0
13 Logic Switch~
5 152 164 0 1 11
0 9
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 A
-4 -19 3 -11
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
43551.5 0
0
13 Logic Switch~
5 152 205 0 1 11
0 8
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 B
-9 -18 -2 -10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3124 0 0
2
43551.5 0
0
14 Logic Display~
6 765 298 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
7 CarryOu
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3421 0 0
2
43551.5 0
0
14 Logic Display~
6 628 213 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
6 SumOut
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
43551.5 0
0
5 4081~
219 522 314 0 3 22
0 7 6 4
0
0 0 624 0
4 4081
-7 -24 21 -16
4 AndB
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
5572 0 0
2
43551.5 0
0
5 4081~
219 364 302 0 3 22
0 9 8 5
0
0 0 624 0
4 4081
-7 -24 21 -16
4 AndA
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
8901 0 0
2
43551.5 0
0
5 4071~
219 656 312 0 3 22
0 4 5 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
7361 0 0
2
43551.5 0
0
5 4030~
219 516 233 0 3 22
0 7 6 3
0
0 0 624 0
4 4030
-7 -24 21 -16
4 XorB
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
4747 0 0
2
43551.5 0
0
5 4030~
219 358 196 0 3 22
0 9 8 7
0
0 0 624 0
4 4030
-7 -24 21 -16
4 XorA
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
972 0 0
2
43551.5 0
0
12
3 1 2 0 0 4224 0 8 4 0 0 5
689 312
753 312
753 324
765 324
765 316
3 1 3 0 0 4224 0 9 5 0 0 5
549 233
616 233
616 239
628 239
628 231
3 1 4 0 0 4224 0 6 8 0 0 4
543 314
635 314
635 303
643 303
3 2 5 0 0 16512 0 7 8 0 0 7
385 302
385 345
494 345
494 389
635 389
635 321
643 321
0 2 6 0 0 8192 0 0 6 9 0 3
418 247
418 323
498 323
0 1 7 0 0 4224 0 0 6 10 0 3
461 196
461 305
498 305
0 2 8 0 0 4096 0 0 7 11 0 3
246 205
246 311
340 311
0 1 9 0 0 4096 0 0 7 12 0 3
266 164
266 293
340 293
1 2 6 0 0 4224 0 1 9 0 0 4
161 247
492 247
492 242
500 242
3 1 7 0 0 0 0 10 9 0 0 4
391 196
492 196
492 224
500 224
1 2 8 0 0 4224 0 3 10 0 0 2
164 205
342 205
1 1 9 0 0 4224 0 2 10 0 0 4
164 164
334 164
334 187
342 187
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
