CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
213 80 1278 963
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
381 176 494 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 159 178 0 1 11
0 2
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6748 0 0
2
43551.5 0
0
13 Logic Switch~
5 89 178 0 1 11
0 9
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6901 0 0
2
43551.5 0
0
5 4071~
219 630 258 0 3 22
0 7 6 5
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
842 0 0
2
43551.5 0
0
5 4081~
219 441 367 0 3 22
0 3 2 4
0
0 0 624 0
4 4081
-7 -24 21 -16
4 AndC
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
3277 0 0
2
43551.5 0
0
5 4081~
219 442 268 0 3 22
0 8 9 6
0
0 0 624 0
4 4081
-7 -24 21 -16
4 AndB
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
4212 0 0
2
43551.5 0
0
5 4081~
219 439 175 0 3 22
0 2 3 7
0
0 0 624 0
4 4081
-7 -24 21 -16
4 AndA
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
4720 0 0
2
43551.5 0
0
9 Inverter~
13 278 284 0 2 22
0 2 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NotB
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
5551 0 0
2
43551.5 0
0
9 Inverter~
13 271 218 0 2 22
0 9 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NotA
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
6986 0 0
2
43551.5 0
0
14 Logic Display~
6 547 355 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
6 Borrow
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8745 0 0
2
43551.5 0
0
14 Logic Display~
6 730 241 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
7 DiffOut
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9592 0 0
2
43551.5 0
0
12
0 2 2 0 0 8336 0 0 4 11 0 3
171 283
171 376
417 376
0 1 3 0 0 4224 0 0 4 8 0 3
320 218
320 358
417 358
3 1 4 0 0 4224 0 4 9 0 0 5
462 367
535 367
535 381
547 381
547 373
3 1 5 0 0 4224 0 3 10 0 0 5
663 258
718 258
718 267
730 267
730 259
3 2 6 0 0 4224 0 5 3 0 0 4
463 268
609 268
609 267
617 267
3 1 7 0 0 4224 0 6 3 0 0 4
460 175
542 175
542 249
617 249
0 1 2 0 0 0 0 0 6 11 0 4
171 192
358 192
358 166
415 166
2 2 3 0 0 0 0 8 6 0 0 4
292 218
407 218
407 184
415 184
2 1 8 0 0 4224 0 7 5 0 0 4
299 284
405 284
405 259
418 259
0 2 9 0 0 8192 0 0 5 12 0 5
244 218
244 247
347 247
347 277
418 277
1 1 2 0 0 0 0 1 7 0 0 3
171 178
171 284
263 284
1 1 9 0 0 12416 0 2 8 0 0 4
101 178
102 178
102 218
256 218
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
