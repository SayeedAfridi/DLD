CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 963
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 63 290 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
3 Bin
-16 -18 5 -10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43555.5 0
0
13 Logic Switch~
5 65 243 0 1 11
0 9
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 B
-9 -21 -2 -13
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
391 0 0
2
43555.5 0
0
13 Logic Switch~
5 63 197 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21104 0
2 5V
-6 -16 8 -8
1 A
-10 -18 -3 -10
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3124 0 0
2
43555.5 0
0
14 Logic Display~
6 793 317 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Bout
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3421 0 0
2
43555.5 0
0
14 Logic Display~
6 666 203 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Sout
-14 -21 14 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
43555.5 0
0
9 Inverter~
13 468 319 0 2 22
0 8 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
5572 0 0
2
43555.5 0
0
9 Inverter~
13 218 326 0 2 22
0 11 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
8901 0 0
2
43555.5 0
0
5 4071~
219 689 329 0 3 22
0 4 5 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
7361 0 0
2
43555.5 0
0
5 4081~
219 553 329 0 3 22
0 7 6 4
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
4747 0 0
2
43555.5 0
0
5 4081~
219 318 341 0 3 22
0 10 9 5
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
43555.5 0
0
5 4030~
219 537 221 0 3 22
0 8 6 3
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
3472 0 0
2
43555.5 0
0
5 4030~
219 310 222 0 3 22
0 11 9 8
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
9998 0 0
2
43555.5 0
0
14
3 1 2 0 0 4224 0 8 4 0 0 5
722 329
781 329
781 343
793 343
793 335
3 1 3 0 0 4224 0 11 5 0 0 5
570 221
654 221
654 229
666 229
666 221
3 1 4 0 0 4224 0 9 8 0 0 4
574 329
668 329
668 320
676 320
3 2 5 0 0 8320 0 10 8 0 0 5
339 341
339 374
668 374
668 338
676 338
0 2 6 0 0 8192 0 0 9 8 0 3
390 290
390 338
529 338
2 1 7 0 0 4224 0 6 9 0 0 4
489 319
521 319
521 320
529 320
0 1 8 0 0 4096 0 0 6 9 0 3
429 222
429 319
453 319
1 2 6 0 0 4224 0 1 11 0 0 4
75 290
513 290
513 230
521 230
3 1 8 0 0 4224 0 12 11 0 0 4
343 222
513 222
513 212
521 212
0 2 9 0 0 8192 0 0 10 13 0 3
117 243
117 350
294 350
2 1 10 0 0 4224 0 7 10 0 0 4
239 326
286 326
286 332
294 332
0 1 11 0 0 4096 0 0 7 14 0 3
165 197
165 326
203 326
1 2 9 0 0 4224 0 2 12 0 0 4
77 243
286 243
286 231
294 231
1 1 11 0 0 4224 0 3 12 0 0 4
75 197
286 197
286 213
294 213
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
