CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 963
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 342 192 0 1 11
0 4
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
317 0 0
2
43551.5 0
0
13 Logic Switch~
5 266 192 0 1 11
0 5
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3108 0 0
2
43551.5 0
0
14 Logic Display~
6 714 384 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
7 CArryOu
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4299 0 0
2
43551.5 0
0
14 Logic Display~
6 876 277 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
6 SumOut
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9672 0 0
2
43551.5 0
0
5 4071~
219 721 300 0 3 22
0 3 2 9
0
0 0 624 0
4 4071
-7 -24 21 -16
3 OrA
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
7876 0 0
2
43551.5 0
0
5 4081~
219 556 396 0 3 22
0 5 4 8
0
0 0 624 0
4 4081
-7 -24 21 -16
4 AndC
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
6369 0 0
2
43551.5 0
0
5 4081~
219 551 309 0 3 22
0 5 6 2
0
0 0 624 0
4 4081
-7 -24 21 -16
4 AndB
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
9172 0 0
2
43551.5 0
0
5 4081~
219 550 217 0 3 22
0 7 4 3
0
0 0 624 0
4 4081
-7 -24 21 -16
4 AndA
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
7100 0 0
2
43551.5 0
0
9 Inverter~
13 413 273 0 2 22
0 4 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NotB
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
3820 0 0
2
43551.5 0
0
9 Inverter~
13 412 218 0 2 22
0 5 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
4 NotA
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7678 0 0
2
43551.5 0
0
12
3 2 2 0 0 4224 0 7 5 0 0 2
572 309
708 309
3 1 3 0 0 12432 0 8 5 0 0 4
571 217
579 217
579 291
708 291
2 0 4 0 0 4224 0 6 0 0 10 3
532 405
354 405
354 272
0 1 5 0 0 8320 0 0 6 6 0 3
277 300
277 387
532 387
2 2 6 0 0 12416 0 9 7 0 0 4
434 273
435 273
435 318
527 318
0 1 5 0 0 0 0 0 7 9 0 3
277 218
277 300
527 300
0 2 4 0 0 0 0 0 8 10 0 4
354 232
518 232
518 226
526 226
2 1 7 0 0 4224 0 10 8 0 0 4
433 218
518 218
518 208
526 208
1 1 5 0 0 0 0 2 10 0 0 4
278 192
277 192
277 218
397 218
1 1 4 0 0 0 0 1 9 0 0 3
354 192
354 273
398 273
3 1 8 0 0 4224 0 6 3 0 0 5
577 396
702 396
702 410
714 410
714 402
3 1 9 0 0 4224 0 5 4 0 0 3
754 300
876 300
876 295
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
