CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1278 963
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 194 270 0 1 11
0 7
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3171 0 0
2
43551.5 0
0
13 Logic Switch~
5 193 211 0 1 11
0 8
0
0 0 21104 0
2 0V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4139 0 0
2
43551.5 0
0
14 Logic Display~
6 952 305 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
7 BorrowO
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6435 0 0
2
43551.5 0
0
14 Logic Display~
6 942 166 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
7 Differe
-24 -21 25 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5283 0 0
2
43551.5 0
0
5 4011~
219 721 187 0 3 22
0 5 4 3
0
0 0 624 0
4 4011
-7 -24 21 -16
5 And1A
-18 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
6874 0 0
2
43551.5 0
0
5 4011~
219 790 310 0 3 22
0 4 4 2
0
0 0 624 0
4 4011
-7 -24 21 -16
4 AndD
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 4 1 0
1 U
5305 0 0
2
43551.5 1
0
5 4011~
219 494 161 0 3 22
0 8 6 5
0
0 0 624 0
4 4011
-7 -24 21 -16
4 AndC
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 3 1 0
1 U
34 0 0
2
43551.5 0
0
5 4011~
219 496 308 0 3 22
0 6 7 4
0
0 0 624 0
4 4011
-7 -24 21 -16
4 AndB
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 1 0
1 U
969 0 0
2
43551.5 0
0
5 4011~
219 346 247 0 3 22
0 8 7 6
0
0 0 624 0
4 4011
-7 -24 21 -16
4 AndA
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 1 0
1 U
8402 0 0
2
43551.5 0
0
12
3 1 2 0 0 4224 0 6 3 0 0 5
817 310
940 310
940 331
952 331
952 323
3 1 3 0 0 4224 0 5 4 0 0 3
748 187
942 187
942 184
0 0 4 0 0 8192 0 0 0 4 5 3
689 308
689 307
758 307
3 2 4 0 0 4224 0 8 5 0 0 4
523 308
689 308
689 196
697 196
2 1 4 0 0 0 0 6 6 0 0 4
766 319
758 319
758 301
766 301
3 1 5 0 0 4224 0 7 5 0 0 4
521 161
689 161
689 178
697 178
3 0 6 0 0 4096 0 9 0 0 8 2
373 247
462 247
1 2 6 0 0 8320 0 8 7 0 0 4
472 299
462 299
462 170
470 170
0 2 7 0 0 8320 0 0 8 11 0 3
274 270
274 317
472 317
0 1 8 0 0 8320 0 0 7 12 0 3
291 211
291 152
470 152
1 2 7 0 0 0 0 1 9 0 0 4
206 270
314 270
314 256
322 256
1 1 8 0 0 0 0 2 9 0 0 4
205 211
314 211
314 238
322 238
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
